`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:47:05 05/09/2014 
// Design Name: 
// Module Name:    lp 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ring_counter(
input clk,
input reset,
output  [1:0] selector 
    );
//wire [1:0] counter_out;
//UpCounter_SyncReset two_bit_counter(clk,reset,selector);
//dec2x4 rotating (counter_out,selector);
endmodule
